//~ `New testbench
`timescale  1ns / 1ps

module tb_CNN;

// CNN Parameters
parameter PERIOD  = 10;


// CNN Inputs
reg   clk                                  = 0 ;
reg   rstn                                 = 0 ;
reg   [44:0]  weight_m_1                   = {9'd2,9'd5,9'd4,9'd5,9'd6} ;
reg   [44:0]  weight_m_2                   = {9'd3,9'd3,9'd2,9'd5,9'd6} ;
reg   [44:0]  weight_m_3                   = {9'd5,9'd3,9'd3,9'd2,9'd6} ;
reg   [44:0]  weight_m_4                   = {9'd4,9'd1,9'd1,9'd5,9'd3} ;
reg   [44:0]  weight_m_5                   = {9'd2,9'd3,9'd8,9'd5,9'd1} ;
reg   signed [8:0]  bias                          = 9'd38 ;

// CNN Outputs
wire  conv_valid                                 ;
wire  signed [21:0]  conv_data                   ;

initial
begin
    forever #(PERIOD/2)  clk=~clk;
end

initial
begin
    #(PERIOD*2) rstn  =  1;
end

 // 定义一个5x5x6的三维数组
    reg signed [8:0] conv1_weight [0:4][0:4][0:5]; 
    reg signed [44:0] conv1_weight_1_m_n [0:4];

    parameter filename = "E:/spyder/matlab/conv1_weight_data.txt";
    integer fid; // 文件句柄
    integer i,j,k; // 
    initial begin
        fid = $fopen(filename, "r");
        
            if(fid != 0) begin
                for(i=0;i<6;i = i + 1) begin
                    for (j = 0; j<5; j = j + 1) begin
                        for (k = 0; k<5; k = k + 1) begin
                            $fscanf(fid, "%b\n", conv1_weight[j][k][i]);
                        end

                    end
                end
            end 

        $fclose(fid);

    end

    initial begin
        #30
            for (j = 0; j<5; j = j + 1) begin
                for (k = 0; k<5; k = k + 1) begin
                    // #1
                    conv1_weight_1_m_n[j] = {conv1_weight_1_m_n[j][35:0],conv1_weight[k][j][0]};
                end
                
            end
    end


CNN  u_CNN (
    .clk                     ( clk                ),
    .rstn                    ( rstn               ),
    .weight_m_1              ( weight_m_1  [44:0] ),
    .weight_m_2              ( weight_m_2  [44:0] ),
    .weight_m_3              ( weight_m_3  [44:0] ),
    .weight_m_4              ( weight_m_4  [44:0] ),
    .weight_m_5              ( weight_m_5  [44:0] ),
    .bias                    ( bias        [8:0]  ),
    .conv_valid              ( conv_valid         ),
    .conv_data               ( conv_data          )
);

always @(*) begin
    weight_m_1 <= conv1_weight_1_m_n[0];
    weight_m_2 <= conv1_weight_1_m_n[1];
    weight_m_3 <= conv1_weight_1_m_n[2];
    weight_m_4 <= conv1_weight_1_m_n[3];
    weight_m_5 <= conv1_weight_1_m_n[4];
end

    integer file_conv1;
    initial begin
        #10
        file_conv1 = $fopen("E:/spyder/FPGA/src/TXT/conv1_data_check.txt","w");
    end

    reg [9:0] conv_data_cnt;
    reg write_flag;
    always @(posedge clk or negedge rstn) begin
        if(rstn == 1'b0) begin
                conv_data_cnt<= 0;
                write_flag <= 1;
            end
        else if(conv_valid&&write_flag) begin 
                $fwrite(file_conv1, "%-15d\n", conv_data);
                conv_data_cnt <= conv_data_cnt + 1;
            end
        else if(conv_data_cnt == 28*28) begin
                conv_data_cnt<= 0;
                write_flag <= 0;
                $fclose(fid);
            end
        else begin
                conv_data_cnt<= conv_data_cnt;
                write_flag <= write_flag;
            end
    end



endmodule